/home/ecegrid/a/mg71/ece337/Lab2/source/tb_adder_nbit.sv