/home/ecegrid/a/mg71/ece337/Lab2/source/adder_1bit.sv