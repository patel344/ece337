// $Id: $
// File name:   sensor_d.sv
// Created:     1/17/2017
// Author:      Parth Patel
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: Dataflow Style Sensor Error Detector.
