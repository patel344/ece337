// $Id: $
// File name:   sensor_s.sv
// Created:     1/17/2017
// Author:      Parth Patel
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: Structural Style Sensor Error Detector module.
